-- assembled from test_prog.asm on 2015-04-16 11:45:07.910319 CEST

--  Address    Code        Basic                     Source
-- 
-- 0x00000000  0x340200c8  ori $2,$0,0x000000c8  6         ori $2,$0, 200  # set eight registers for test purpose, do not use $0 and $1
-- 0x00000004  0x34030032  ori $3,$0,0x00000032  7         ori $3,$0, 50
-- 0x00000008  0x340403ff  ori $4,$0,0x000003ff  8         ori $4,$0, 1023 # stores add result (2000 + 50)
-- 0x0000000c  0x340503ff  ori $5,$0,0x000003ff  9         ori $5,$0, 1023 # stores addi result(2000 + 2000 ie)
-- 0x00000010  0x340603ff  ori $6,$0,0x000003ff  10        ori $6,$0, 1023 # stores divu result(2000 / 50)
-- 0x00000014  0x340703ff  ori $7,$0,0x000003ff  11        ori $7,$0, 1023 # stores mult result(2000 * 50)
-- 0x00000018  0x340803ff  ori $8,$0,0x000003ff  12        ori $8,$0, 1023 # stores sub result(2000 - 50)
-- 0x0000001c  0x34090076  ori $9,$0,0x00000076  15        ori $9,$0, 118   # ( 0b01110110 ) 
-- 0x00000020  0x340a00b0  ori $10,$0,0x000000b0 16        ori $10,$0, 176  # ( 0b10101010 )
-- 0x00000024  0x340b03ff  ori $11,$0,0x000003ff 17        ori $11,$0, 1023 # stores and result (118 & 176)
-- 0x00000028  0x340c03ff  ori $12,$0,0x000003ff 18        ori $12,$0, 1023 # stores andi result(118 & 225 ie)
-- 0x0000002c  0x340d03ff  ori $13,$0,0x000003ff 19        ori $13,$0, 1023 # stores or result()
-- 0x00000030  0x340d03ff  ori $13,$0,0x000003ff 21        ori $13,$0, 1023 # stores arithmetic branch condition
-- 0x00000034  0x340d03ff  ori $13,$0,0x000003ff 22        ori $13,$0, 1023 # stores logic branch condition
-- 0x00000038  0x201403fc  addi $20,$0,0x000003fc26        addi $20, $0, 1020    # .data offset voor "hardware"
-- 0x0000003c  0xae82ffe8  sw $2,0xffffffe8($20) 28        sw   $2, -24($20) # store all the registers to the memory, offset and register flipped in order to switch easy between simulator and hardware
-- 0x00000040  0xae83ffec  sw $3,0xffffffec($20) 29        sw   $3, -20($20)
-- 0x00000044  0xae84fff0  sw $4,0xfffffff0($20) 30        sw   $4, -16($20)
-- 0x00000048  0xae85fff4  sw $5,0xfffffff4($20) 31        sw   $5, -12($20)
-- 0x0000004c  0xae86fff8  sw $6,0xfffffff8($20) 32        sw   $6, -8($20)
-- 0x00000050  0xae87fffc  sw $7,0xfffffffc($20) 33        sw   $7, -4($20)
-- 0x00000054  0xae880000  sw $8,0x00000000($20) 34        sw   $8, 0($20)
-- 0x00000058  0x8e82ffe8  lw $2,0xffffffe8($20) 37        lw   $2, -24($20) # load all the register from the memory
-- 0x0000005c  0x8e83ffec  lw $3,0xffffffec($20) 38        lw   $3, -20($20)
-- 0x00000060  0x8e84fff0  lw $4,0xfffffff0($20) 39        lw   $4, -16($20)
-- 0x00000064  0x8e85fff4  lw $5,0xfffffff4($20) 40        lw   $5, -12($20)
-- 0x00000068  0x8e86fff8  lw $6,0xfffffff8($20) 41        lw   $6, -8($20)
-- 0x0000006c  0x8e87fffc  lw $7,0xfffffffc($20) 42        lw   $7, -4($20)
-- 0x00000070  0x8e880000  lw $8,0x00000000($20) 43        lw   $8, 0($20) 
-- 0x00000074  0x00432020  add $4,$2,$3          45        add    $4, $2, $3  
-- 0x00000078  0x20a60032  addi $6,$5,0x00000032 46        addi   $6, $5, 50
-- 0x0000007c  0x00c74024  and $8,$6,$7          48        and    $8, $6, $7
-- 0x00000080  0x3043aaaa  andi $3,$2,0x0000aaaa 49        andi   $3, $2, 0xAAAA
-- 0x00000084  0x10640001  beq $3,$4,0x00000001  51        beq    $3, $4, branch1 ## 
-- 0x00000088  0x10640000  beq $3,$4,0x00000000  52        beq    $3, $4, branch1 ## 
-- 0x0000008c  0x1cc00001  bgtz $6,0x00000001    54        bgtz   $6, branch2
-- 0x00000090  0x1cc00000  bgtz $6,0x00000000    55        bgtz   $6, branch2     ## duplicat both to verify right behaviour
-- 0x00000094  0x0107001b  divu $8,$7            58        divu   $8, $7
-- 0x00000098  0x00003810  mfhi $7               59        mfhi   $7
-- 0x0000009c  0x00004012  mflo $8               60        mflo   $8
-- 0x000000a0  0x00430018  mult $2,$3            63        mult   $2, $3
-- 0x000000a4  0x00001010  mfhi $2               64        mfhi   $2
-- 0x000000a8  0x00001812  mflo $3               65        mflo   $3
-- 0x000000ac  0x00000000  nop                   67        nop	   	
-- 0x000000b0  0x00000000  nop                   68        nop	
-- 0x000000b4  0xae82ffe8  sw $2,0xffffffe8($20) 70        sw   $2, -24($20)
-- 0x000000b8  0xae83ffec  sw $3,0xffffffec($20) 71        sw   $3, -20($20)
-- 0x000000bc  0xae84fff0  sw $4,0xfffffff0($20) 72        sw   $4, -16($20)
-- 0x000000c0  0xae85fff4  sw $5,0xfffffff4($20) 73        sw   $5, -12($20)
-- 0x000000c4  0xae86fff8  sw $6,0xfffffff8($20) 74        sw   $6, -8($20)
-- 0x000000c8  0xae87fffc  sw $7,0xfffffffc($20) 75        sw   $7, -4($20)
-- 0x000000cc  0xae880000  sw $8,0x00000000($20) 76        sw   $8, 0($20) # load some registers
-- 0x000000d0  0x08000016  j 0x00000058          81        j begin ## jump to start
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
PACKAGE program IS
	CONSTANT low_address	: INTEGER := 0; 
	CONSTANT high_address	: INTEGER := 255;

	TYPE mem_array IS ARRAY (low_address TO high_address) OF std_logic_vector(31 DOWNTO 0);
	CONSTANT program : mem_array := (
"00110100000000100000000011001000",
"00110100000000110000000000110010",
"00110100000001000000001111111111",
"00110100000001010000001111111111",
"00110100000001100000001111111111",
"00110100000001110000001111111111",
"00110100000010000000001111111111",
"00110100000010010000000001110110",
"00110100000010100000000010110000",
"00110100000010110000001111111111",
"00110100000011000000001111111111",
"00110100000011010000001111111111",
"00110100000011010000001111111111",
"00110100000011010000001111111111",
"00100000000101000000001111111100",
"10101110100000101111111111101000",
"10101110100000111111111111101100",
"10101110100001001111111111110000",
"10101110100001011111111111110100",
"10101110100001101111111111111000",
"10101110100001111111111111111100",
"10101110100010000000000000000000",
"10001110100000101111111111101000",
"10001110100000111111111111101100",
"10001110100001001111111111110000",
"10001110100001011111111111110100",
"10001110100001101111111111111000",
"10001110100001111111111111111100",
"10001110100010000000000000000000",
"00000000010000110010000000100000",
"00100000101001100000000000110010",
"00000000110001110100000000100100",
"00110000010000111010101010101010",
"00010000011001000000000000000001",
"00010000011001000000000000000000",
"00011100110000000000000000000001",
"00011100110000000000000000000000",
"00000001000001110000000000011011",
"00000000000000000011100000010000",
"00000000000000000100000000010010",
"00000000010000110000000000011000",
"00000000000000000001000000010000",
"00000000000000000001100000010010",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"10101110100000101111111111101000",
"10101110100000111111111111101100",
"10101110100001001111111111110000",
"10101110100001011111111111110100",
"10101110100001101111111111111000",
"10101110100001111111111111111100",
"10101110100010000000000000000000",
"00001000000000000000000000010110",

OTHERS => "00000000000000000000000000000000");

END;
