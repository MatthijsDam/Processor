--------------------------------------------------------------
-- 
-- Clock driven Memory (results in 1 clockcycle delay) 
--
--------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.ALL;

ENTITY memory IS
	PORT(
		address_bus	: IN  std_logic_vector(31 DOWNTO 0);
		databus_in	: IN  std_logic_vector(31 DOWNTO 0);
		databus_out : OUT std_logic_vector(31 DOWNTO 0);
		write		: IN  std_logic;
		clk			: IN  std_logic
	);
END memory;

ARCHITECTURE behaviour OF memory IS
	CONSTANT low_address	: INTEGER := 0; 
	CONSTANT high_address	: INTEGER := 255;

	TYPE mem_array IS ARRAY (low_address TO high_address) OF std_logic_vector(31 DOWNTO 0);
	
	SIGNAL mem 		: mem_array := 
					 ("00110100000000100000011111010000",
						"00110100000000110000000000110010",
						"00110100000010010000000001110110",
						"00110100000010100000000010110000",
						"00110100000011100000000000000000",
						"00110100000011110000000000000000",
						"00110100000100000000000000000001",
						"00110100000110100000000000000000",
						"00110100000110110000000000000000",
						"00100000000101000000001111111100",
						"10101110100000100000000000000000",
						"10101110100000111111111111111100",
						"10101110100010011111111111100100",
						"10101110100010101111111111100000",
						"10001110100000100000000000000000",
						"10001110100000111111111111111100",
						"00000000010000110010000000100000",
						"00100000010001010000011111010000",
						"00000000011000100000000000011011",
						"00000000000000000011000000010000",
						"00000000010000110000000000011000",
						"00000000000000000011100000010010",
						"00000000010000110100000000100010",
						"00100011010110100000000000000001",
						"00000001110100000111000000100110",
						"10101110100001001111111111111000",
						"10101110100001011111111111110100",
						"10101110100001101111111111110000",
						"10101110100001111111111111101100",
						"10101110100010001111111111101000",
						"10101110100110101111111111010000",
						"00010001110000001111111111101110",
						"10001110100010011111111111100100",
						"10001110100010101111111111100000",
						"00000001001010100101100000100100",
						"00110001001011000000000010110111",
						"00000001001010100110100000100101",
						"00100011011110110000000000000001",
						"00000001111100000111100000100110",
						"10101110100010111111111111011100",
						"10101110100011001111111111011000",
						"10101110100011011111111111010100",
						"10101110100110111111111111001100",
						"00011101111000001111111111110100",
						"00001000000000000000000000001110",
						OTHERS => "00000000000000000000000000000000"
						);

	
	BEGIN
		PROCESS(clk,address_bus)
			VARIABLE address 	: INTEGER;
	
		BEGIN
			IF to_integer(unsigned(address_bus(31 DOWNTO 2))) <= high_address THEN
				address 	:=  to_integer(unsigned(address_bus(31 DOWNTO 2)));
			END	IF;
			databus_out <= mem(address);
			IF rising_edge(clk) THEN
				IF write = '1' THEN
					mem(address) <= databus_in;			
				END IF;
			END IF;
		END PROCESS;

END ARCHITECTURE;


