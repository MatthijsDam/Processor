--------------------------------------------------------------
-- 
-- Clock driven Memory (results in 1 clockcycle delay) 
--
--------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.ALL;

ENTITY memory IS
	PORT(
		address_bus	: IN  std_logic_vector(31 DOWNTO 0);
		databus_in	: IN  std_logic_vector(31 DOWNTO 0);
		databus_out : OUT std_logic_vector(31 DOWNTO 0);
		write		: IN  std_logic;
		clk			: IN  std_logic
	);
END memory;

ARCHITECTURE behaviour OF memory IS
	CONSTANT low_address	: INTEGER := 0; 
	CONSTANT high_address	: INTEGER := 256;

	TYPE mem_array IS ARRAY (low_address TO high_address) OF std_logic_vector(31 DOWNTO 0);
	
	SIGNAL mem 		: mem_array := 
					 ("00110100000000100000000011001000",
						"00110100000000110000000000110010",
						"00110100000001000000001111111111",
						"00110100000001010000001111111111",
						"00110100000001100000001111111111",
						"00110100000001110000001111111111",
						"00110100000010000000001111111111",
						"00110100000010010000000001110110",
						"00110100000010100000000010110000",
						"00110100000010110000001111111111",
						"00110100000011000000001111111111",
						"00110100000011010000001111111111",
						"00110100000011010000001111111111",
						"00110100000011010000001111111111",
						"00100000000101000000000100000000",
						"10101110100000101111111111101000",
						"10101110100000111111111111101100",
						"10101110100001001111111111110000",
						"10101110100001011111111111110100",
						"10101110100001101111111111111000",
						"10101110100001111111111111111100",
						"10101110100010000000000000000000",
						"10001110100000101111111111101000",
						"10001110100000111111111111101100",
						"10001110100001001111111111110000",
						"10001110100001011111111111110100",
						"10001110100001101111111111111000",
						"10001110100001111111111111111100",
						"10001110100010000000000000000000",
						"00000000010000110010000000100000",
						"00100000101001100000000000110010",
						"00000000110001110100000000100100",
						"00110000010000111010101010101010",
						"00010000011001000000000000000001",
						"00010000011001000000000000000000",
						"00011100110000000000000000000001",
						"00011100110000000000000000000000",
						"00000001000001110000000000011011",
						"00000000000000000011100000010000",
						"00000000000000000100000000010010",
						"00000000010000110000000000011000",
						"00000000000000000001000000010000",
						"00000000000000000001100000010010",
						"00000000000000000000000000000000",
						"00000000000000000000000000000000",
						"10101110100000101111111111101000",
						"10101110100000111111111111101100",
						"10101110100001001111111111110000",
						"10101110100001011111111111110100",
						"10101110100001101111111111111000",
						"10101110100001111111111111111100",
						"10101110100010000000000000000000",
						"00001000000100000000000000010110",
					  OTHERS => "00000000000000000000000000000000"
						);

	
	BEGIN
		PROCESS(clk,address_bus)
			VARIABLE address 	: INTEGER;
	
		BEGIN
			IF to_integer(unsigned(address_bus(31 DOWNTO 2))) < high_address THEN
				address 	:=  to_integer(unsigned(address_bus(31 DOWNTO 2)));
			END	IF;
			databus_out <= mem(address);
			IF rising_edge(clk) THEN
				IF write = '1' THEN
					mem(address) <= databus_in;			
				END IF;
			END IF;
		END PROCESS;

END ARCHITECTURE;


