--------------------------------------------------------------
-- 
-- Processor
--
--------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE work.ALL;
USE intruction_decode_defs.ALL;


ENTITY processor IS
    PORT(
        address_bus     : OUT std_logic_vector(31 DOWNTO 0);
        databus_in      : IN  std_logic_vector(31 DOWNTO 0);
        databus_out     : OUT std_logic_vector(31 DOWNTO 0);
        read            : OUT std_logic;
        write           : OUT std_logic;
        reset           : IN  std_logic;
        clk             : IN  std_logic
    );
END processor;

ARCHITECTURE behaviour OF processor IS
    TYPE fsm_state_t IS (fetch, execute, mem);
    TYPE reg_bank_t IS ARRAY (0 TO 31) OF std_logic_vector(31 DOWNTO 0); 
    SIGNAL reg                      : reg_bank_t := 
         ("00000000000000000000000000000000",
          "00000000000000000000000000000001",
          "00000000000000000000000000000010",
          OTHERS => "00000000000000000000000000000000"
          );
          
    SIGNAL reg_LO, reg_HI     : std_logic_vector(31 DOWNTO 0);
      SIGNAL state              : fsm_state_t;
    
BEGIN


    PROCESS(clk,reset)
        VARIABLE pc                 : INTEGER := 0;
        VARIABLE instruction        : std_logic_vector(31 DOWNTO 0);
       
        VARIABLE opcode             : std_logic_vector(5 DOWNTO 0);

        VARIABLE src                : INTEGER RANGE 0 TO 31;
        VARIABLE src_tgt            : INTEGER RANGE 0 TO 31;
        VARIABLE dst                : INTEGER RANGE 0 TO 31;
        
        VARIABLE operand1           : std_logic_vector(31 DOWNTO 0);
        VARIABLE operand2           : std_logic_vector(31 DOWNTO 0);
        
        VARIABLE funct              : std_logic_vector(5 DOWNTO 0);

        VARIABLE imm                : std_logic_vector(15 DOWNTO 0);
        VARIABLE target             : std_logic_vector(25 DOWNTO 0);
        VARIABLE temp64             : std_logic_vector(63 DOWNTO 0);

        

    -- A read operation has 1 clock cycle delay
    PROCEDURE memory_read(
                pc      : IN INTEGER; 
                data    : OUT std_logic_vector(31 DOWNTO 0)) IS
        
        VARIABLE address     : std_logic_vector(31 DOWNTO 0);

        BEGIN
            read        <= '1';
            address     := std_logic_vector(to_unsigned(pc,30)) & "00";
            address_bus <= address;
            data        := databus_in;
    END memory_read;

    PROCEDURE memory_write(
                    address : IN std_logic_vector(31 DOWNTO 0); 
                    data    : IN std_logic_vector(31 DOWNTO 0)) IS    
        BEGIN
            write         <= '1';
            databus_out <= data;
    END memory_write;  
      

    BEGIN
        IF reset='1' THEN 
            state           <= fetch;
            pc              := 0;
            read            <= '0';
            write           <= '0';
            databus_out     <= "UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU";
            address_bus     <= "UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU";


            
        ELSIF rising_edge(clk) THEN
            CASE state IS
                WHEN fetch =>
                    --
                    -- Instruction fetch
                    --
                    memory_read(pc,instruction);

                    -- Increase program counter
                    pc := pc+1;

                    state <= execute;

                WHEN execute =>
                    state <= fetch; ---- let op!
                  
                    -- Common
                    opcode      := instruction(31 DOWNTO 26);

                    -- Common R and I
                    src         := to_integer(unsigned(instruction(25 DOWNTO 21)));
                    src_tgt     := to_integer(unsigned(instruction(20 DOWNTO 16)));
                    
                    -- Both registers (R-Type):
                    dst         := to_integer(unsigned(instruction(15 DOWNTO 11)));
                    funct       := instruction( 5 DOWNTO  0);
                    -----------------------------------------
                    -- One immediate (I-Type):
                    imm         := std_logic_vector(resize(signed(instruction(15 DOWNTO 0)),32));
                    -----------------------------------------
                    -- Jump (J-Type):
                    target      := instruction(25 DOWNTO 0);
                    -----------------------------------------
                    
                    -- Decoding and execution
                    CASE opcode IS
                     -- Arithmetic registers operation or nop
                     WHEN Rtype =>
                        operand1 := reg(src);
                        operand2 := reg(src_tgt);
                       
                        CASE funct IS
                            -- Arithmetic ADD
                            WHEN F_add =>
                                reg(dst) <= std_logic_vector( signed(operand1) + signed(operand2) ); 
                            -- Arithmetic DIVU
                            WHEN F_divu =>
                                --reg(dst) = std_logic_vector( to_unsigned(reg(src), 32) / to_unsigned(reg(src_tgt), 32) ); -- int to logic vector logic needs to be addeda
                            -- Arithmetic MULT
                            WHEN F_mult =>
                                 temp64 := std_logic_vector( signed(operand1) * signed(operand2) ); 
                                 reg_HI <= temp64(63 DOWNTO 32); 
                                 reg_LO <= temp64(31 DOWNTO 0);
                            -- Arithmetic SUB
                            WHEN F_sub =>
                                 reg(dst) <= std_logic_vector( signed(operand1) - signed(operand2) );                                 

                            -- Logic AND
                            WHEN F_and =>      
                                 reg(dst) <= operand1 AND operand2;                                      
                            -- Logic OR
                            WHEN F_or =>
                                 reg(dst) <= operand1 OR operand2 );                                 
                            -- Logic XOR
                            WHEN F_xor =>
                                 reg(dst) <= operand1 XOR operand2 );                                 
                            -- NOP "operation"
                            WHEN F_xor =>
                               --something with reg(0)

                            -- MFHI move from $HI to dst register
                            WHEN F_mfhi =>
                                  reg(dst) <= reg_HI;
                            -- MFLO move from $LO to dst register
                            WHEN F_mflo => 
                                  reg(dst) <= reg_LO;
                            WHEN OTHERS =>     
                        END CASE;

                     -- ADD immediate operation
                     WHEN "001000" =>

                        --reg(src_tgt) = std_logic_vector(reg(src) + imm; -- int to logic vector logic needs to be added
                     -- AND immediate operation
                     WHEN "001100" =>
                        reg(dst) <= operand1(15 DOWNTO 0) AND std_logic_vector(resize(signed(imm),32));
                     -- OR immediate operation
                     WHEN "001101" =>   
                        
                     -- JUMP immediate operation
                     WHEN "000010" =>
                     -- BEQ immediate operation
                     WHEN "000100" =>   
                     -- BGEZ immediate operation
                     WHEN "000001" =>
                     

                     -- LUI immediate operation 
                     WHEN "001111" => 
                        reg(
                     -- Load word  LW memory immediate operation
                     WHEN "100011" =>
                        state <= mem;
                     -- Store word SW memory immediate operation
                     WHEN "101011" => 
                        state <= mem;
                     WHEN OTHERS =>     
                    END CASE;
                WHEN mem =>
                    state <= fetch;
                    
            END CASE;
        END IF;
    END PROCESS;

END ARCHITECTURE;


